interface inter(input logic clk,rst);
  logic [5:0]a;
  logic [5:0]b;
  logic [5:0]y;
  logic sel;
  
endinterface